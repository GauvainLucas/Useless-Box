library verilog;
use verilog.vl_types.all;
entity Servo_vlg_check_tst is
    port(
        PWM             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Servo_vlg_check_tst;
