library verilog;
use verilog.vl_types.all;
entity Bargraph_vlg_vec_tst is
end Bargraph_vlg_vec_tst;
