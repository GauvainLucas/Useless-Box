library verilog;
use verilog.vl_types.all;
entity Servo_vlg_vec_tst is
end Servo_vlg_vec_tst;
